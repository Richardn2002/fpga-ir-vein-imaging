PACKAGE constants IS
    CONSTANT INPUT_X : NATURAL := 128;
    CONSTANT INPUT_Y : NATURAL := 128;

    CONSTANT CLAHE_CLIP_LIMIT : NATURAL := 10;
    CONSTANT CLAHE_PATCH_X_NUM : NATURAL := 4;
    CONSTANT CLAHE_PATCH_Y_NUM : NATURAL := 4;
    CONSTANT CLAHE_PATCH_X : NATURAL := 32;
    CONSTANT CLAHE_PATCH_Y : NATURAL := 32;

    CONSTANT CLAHE_PATCH_ADDR_BITS : NATURAL := 10;
    CONSTANT CLAHE_MAPPING_ADDR_BITS : NATURAL := 8;
    CONSTANT CLAHE_IMG_ADDR_BITS : NATURAL := 14;
    CONSTANT CLAHE_OUTPUT_ADDR_BITS : NATURAL := 14;

    CONSTANT HESSIAN_INPUT_X : NATURAL := (CLAHE_PATCH_X_NUM - 1) * CLAHE_PATCH_X;
    CONSTANT HESSIAN_INPUT_Y : NATURAL := (CLAHE_PATCH_Y_NUM - 1) * CLAHE_PATCH_Y;
    CONSTANT HESSIAN_RADIUS : NATURAL := 3;
    CONSTANT HESSIAN_OUTPUT_X : NATURAL := HESSIAN_INPUT_X - 2 * HESSIAN_RADIUS;
    CONSTANT HESSIAN_OUTPUT_Y : NATURAL := HESSIAN_INPUT_Y - 2 * HESSIAN_RADIUS;
END PACKAGE constants;